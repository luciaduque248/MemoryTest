library verilog;
use verilog.vl_types.all;
entity MemoryTest_vlg_vec_tst is
end MemoryTest_vlg_vec_tst;
