library verilog;
use verilog.vl_types.all;
entity memory_vlg_vec_tst is
end memory_vlg_vec_tst;
