library verilog;
use verilog.vl_types.all;
entity outputPorts_vlg_vec_tst is
end outputPorts_vlg_vec_tst;
